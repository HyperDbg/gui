module sys
fn main() {
	println('hello,world')
}